module sevensegmentsdecoder(
  input logic [3:0] inp,
  output logic [6:0] y
);


always_comb
  begin
  case(inp)
    //                     .abc_defg  
    4'b0000 : y = ~(7'b011_1111);
    4'b0001 : y = ~(7'b000_0110);
    4'b0010 : y = ~(7'b101_1011);
    4'b0011 : y = ~(7'b100_1111);
    4'b0100 : y = ~(7'b110_0110);
    4'b0101 : y = ~(7'b110_1101);
    4'b0110 : y = ~(7'b111_1101);
    4'b0111 : y = ~(7'b000_0111);
    4'b1000 : y = ~(7'b111_1111);
    4'b1001 : y = ~(7'b110_0111);
    4'b1010 : y = ~(7'b111_0111);
    4'b1011 : y = ~(7'b111_1100);
    4'b1100 : y = ~(7'b011_1001);
    4'b1101 : y = ~(7'b101_1110);
	 4'b1110 : y = ~(7'b111_1001);
    4'b1111 : y = ~(7'b111_0001);
	 
  endcase
  end


endmodule 